module CPU ();
  Datapath DP();
  Controller CU();
endmodule // CPU
