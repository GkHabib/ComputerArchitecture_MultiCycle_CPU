module Datapath ();

endmodule // Datapath
