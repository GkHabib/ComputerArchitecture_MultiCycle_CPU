module Controller ();
  
endmodule // Controller
